`timescale 1ns / 1ps

module rdbf;
	reg [935:0] inp;
	reg clk;
	reg high;
	integer i;
    wire [1871:0] out;
    reg [1871:0] mesh;
	reg [467:0] contour;
	reg [935:0] inps[0:1];

	// Instantiate the Unit Under Test (UUT)
	twobit_26x18_mesh uut (
		.inp(inp),
		.clk(clk),
		.high(high),
        .out(out)
	);

    integer i, i_east;
    reg [5:0] ind;

    initial begin
        clk = 0;
        forever begin
            #50 clk = ~clk;
        end
    end

    initial begin
        high = 0;
        inps[1] = 936'b111111111111111111111111111111111111111111111111111111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000011110000000000000000111111111111111100000000000000001111000000000000000011111111111111110000000000000000111100000000000000001111111111111111000000000000000011110000000000000000111111111111111100000000000000001111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111111111111111111111111111111111111111111111111111111;
        inps[0] = 936'b111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111100000000000000000000000000000000111111111111111111110000000000000000000000000000000011111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111100000000000000000000001111111111111111111111111111110000000000000000000000111111111111111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111100000000000000000000000000000000000011111111111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        mesh = 0;
        contour = 468'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    end
    integer select = 0;
	always @(posedge clk) begin
	   high = 1;
	   contour = 468'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        inp = inps[select%2];
        #350;
        mesh = out;
        inp = 0;
        for (i = 467 ; i>=0 ; i=i-1 ) begin
              i_east = (i-i%26)+(i-1+26)%26;
            if((mesh[4*i_east]&mesh[4*i_east+1]&mesh[4*i_east+2]&mesh[4*i_east+3])!=(mesh[4*i]&mesh[4*i+1]&mesh[4*i+2]&mesh[4*i+3])) begin
                if((mesh[4*i]&mesh[4*i+1]&mesh[4*i+2]&mesh[4*i+3]) == 0) begin
                    contour[i] = 1'b0;
                end
                else begin
                    contour[i_east] = 1'b0;
                end
            end
        end
        select = select+1;
        #50;
        mesh = 0;
	end
  
endmodule