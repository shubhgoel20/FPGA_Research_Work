`timescale 1ns / 1ps

module pixel_foll_tb;
	reg [935:0] inp;
	reg clk;
	reg high;
	integer i;
    wire [1871:0] out;
    reg [1871:0] mesh;
	reg [467:0] contour;
	reg [935:0] inps[0:1];

	// Instantiate the Unit Under Test (UUT)
	twobit_26x18_mesh uut (
		.inp(inp),
		.clk(clk),
		.high(high),
        .out(out)
	);

    integer i, i_east, i_south ,x,y;
    reg [5:0] ind;

    task searchneighbour;
        input integer i;

        for( ind=0 ; ind<16 ; ind=ind+1) begin
            case(ind/4)
                0 : begin
                    x = (i-26+468)%468;    //N
                end

                1 : begin
                    x = (i-i%26)+(i+1+26)%26;  //E
                end

                2 : begin
                    x = (i+26+468)%468;    //S
                end

                3 : begin
                    x = (i-i%26)+(i-1+26)%26;  //W
                end
            endcase

            case(ind%4)
                0 : begin
                    y = (x-26+468)%468;    //N
                end

                1 : begin
                    y = (x-x%26)+(x+1+26)%26;  //E
                end

                2 : begin
                    y = (x+26+468)%468;    //S
                end

                3 : begin
                    y = (x-x%26)+(x-1+26)%26;  //W
                end
            endcase

            // Now we will have (x,y) as a pair of neighbours of node (i.e. neighbour1 & neighbour2)

            if (contour[x] != 1'b0) begin
                if ((mesh[4*y]&mesh[4*y+1]&mesh[4*y+2]&mesh[4*y+3])>(mesh[4*x]&mesh[4*x+1]&mesh[4*x+2]&mesh[4*x+3])) begin
                    contour[x] = 1'b0;
                    searchneighbour(x);
                end
            end

        end
        
    endtask
    
    initial begin
        clk = 0;
        forever begin
            #50 clk = ~clk;
        end
    end

    initial begin
        high = 0;
        inps[1] = 936'b111111111111111111111111111111111111111111111111111111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000011110000000000000000111111111111111100000000000000001111000000000000000011111111111111110000000000000000111100000000000000001111111111111111000000000000000011110000000000000000111111111111111100000000000000001111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111111111111111111111111111111111111111111111111111111;
        inps[0] = 936'b111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111100000000000000000000000000000000111111111111111111110000000000000000000000000000000011111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111100000000000000000000001111111111111111111111111111110000000000000000000000111111111111111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111100000000000000000000000000000000000011111111111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        mesh = 0;
        contour = 468'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    end
    integer select = 0;
	always @(posedge clk) begin
	   high = 1;
	   contour = 468'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        inp = inps[select%2];
        #350;
        mesh = out;
        inp = 0;
        for (i = 467 ; i>=0 ; i=i-1 ) begin
              i_east = (i-i%26)+(i-1+26)%26;
              i_south = (i-26+468)%468;

            if(contour[i] != 1'b0) begin            // for i_east
                if((mesh[4*i_east]&mesh[4*i_east+1]&mesh[4*i_east+2]&mesh[4*i_east+3])>(mesh[4*i]&mesh[4*i+1]&mesh[4*i+2]&mesh[4*i+3])) begin
                    contour[i] = 1'b0;
                    searchneighbour(i);
                end

                if(contour[i_east] != 1'b0) begin
                    if((mesh[4*i_east]&mesh[4*i_east+1]&mesh[4*i_east+2]&mesh[4*i_east+3]) < (mesh[4*i]&mesh[4*i+1]&mesh[4*i+2]&mesh[4*i+3])) begin
                        contour[i_east] = 1'b0;
                        searchneighbour(i_east);
                    end
                end
            end

            if(contour[i] != 1'b0) begin            // for i_south
                if((mesh[4*i_south]&mesh[4*i_south+1]&mesh[4*i_south+2]&mesh[4*i_south+3]) > (mesh[4*i]&mesh[4*i+1]&mesh[4*i+2]&mesh[4*i+3])) begin
                    contour[i] = 1'b0;
                    searchneighbour(i);
                end

                if(contour[i_south] != 1'b0) begin
                    if((mesh[4*i_south]&mesh[4*i_south+1]&mesh[4*i_south+2]&mesh[4*i_south+3]) < (mesh[4*i]&mesh[4*i+1]&mesh[4*i+2]&mesh[4*i+3])) begin
                        contour[i_south] = 1'b0;
                        searchneighbour(i_south);
                    end
                end
            end
        end
        select = select+1;
        #50;
        mesh = 0;
	end
  
endmodule