`timescale 1ns / 1ps

module pixel_foll_tb;
	reg [935:0] inp;
	reg clk;
	reg high;
    reg algo; //Controls which algorithm to run. Set it to 0 for pixel foll. and to 1 for RDBF
	integer i;
    
	wire [467:0] contour;
	reg [935:0] inps[0:1];

	// Instantiate the Unit Under Test (UUT)
	twobit_26x18_mesh uut (
		.inp(inp),
		.clk(clk),
		.high(high),
        .algo(algo),
        .contour(contour)
	);

    
    
    initial begin
        clk = 0;
        forever begin
            #50 clk = ~clk;
        end
    end

    initial begin
        algo = 1;
        high = 0;
        inps[1] = 936'b111111111111111111111111111111111111111111111111111111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000011110000000000000000111111111111111100000000000000001111000000000000000011111111111111110000000000000000111100000000000000001111111111111111000000000000000011110000000000000000111111111111111100000000000000001111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111111111111111111111111111111111111111111111111111111;
        inps[0] = 936'b111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111100000000000000000000000000000000111111111111111111110000000000000000000000000000000011111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111100000000000000000000001111111111111111111111111111110000000000000000000000111111111111111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111100000000000000000000000000000000000011111111111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    end
    integer select = 0;
	always @(posedge clk) begin
	   high = 1;
       algo = 1;
        inp = inps[select%2];
        #350;
        select = select+1;
        #50;
	end
  
endmodule