`timescale 1ns / 1ps

module combined_tb;
	reg [935:0] inp; //468 two bit pixel values
	reg clk;
	reg high;
    reg [1:0] algo; // algorithm selector
	integer i;
    
	wire [467:0] contour;
	// reg [935:0] inps[0:1];
    reg [1:0] algos[0:2];
	// Instantiate the Unit Under Test (UUT)
	twobit_26x18_mesh uut (
		.inp(inp),
		.clk(clk),
		.high(high),
        .algo(algo),
        .contour(contour)
	);

    
    
    initial begin
        clk = 0;
        forever begin
            #50 clk = ~clk;
        end
    end

    initial begin
        algo = 2'b00;
        algos[0] = 2'b00;
        algos[1] = 2'b01;
        algos[2] = 2'b10;
        high = 0;
        inp = 936'b111111111111111111111111111111111111111111111111111111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000011110000000000000000111111111111111100000000000000001111000000000000000011111111111111110000000000000000111100000000000000001111111111111111000000000000000011110000000000000000111111111111111100000000000000001111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111111111111111111111111111111111111111111111111111111;

//        inps[1] = 936'b111111111111111111111111111111111111111111111111111111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000011110000000000000000111111111111111100000000000000001111000000000000000011111111111111110000000000000000111100000000000000001111111111111111000000000000000011110000000000000000111111111111111100000000000000001111111111110000000011111111111111110000000011111111111111111111000000001111111111111111000000001111111111111111111100000000111111111111111100000000111111111111111111110000000011111111111111110000000011111111111111111111111111111111111111111111111111111111111111;
//        inps[0] = 936'b111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111100000000000000000000000000000000111111111111111111110000000000000000000000000000000011111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111100000000000000000000001111111111111111111111111111110000000000000000000000111111111111111111111111111111000000000011111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111100000000000000000000000000000000000011111111111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    end

    //algo = 00: Pixel Following
	//algo = 01: RDBF
	//algo = 10: Vertex Following


    integer select = 0;
	always @(posedge clk) begin
	    high = 1;
//      inp = inps[select%2];
        algo = algos[select%3];
//      inp = inps[1];
//      #350;
        select = select+1;
//      #50;
	end
  
endmodule